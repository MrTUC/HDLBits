/*
 * This file could be similar to the previous one. But since the tool sets undefined ports to zero it can just be left empty. This is bad designing habit.
 */

module top_module (
    output zero
);// Module body starts after semicolon
    


endmodule
