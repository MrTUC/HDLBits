/*
 * In this module we connect the input port to the output port. This is done with assigning the input signal to the output signal.
 */

module top_module ( input in, output out );
	assign out = in;
endmodule
